module top_module( 
    input [3:0] in,
    output out_and,
    output out_or,
    output out_xor
);
    assign {out_and,out_or,out_xor} = {(in[3] & in[2] & in[1]&in[0]), (in[3]|in[2]|in[1]|in[0]), (in[3]^in[2]^in[1]^in[0])};
    
endmodule
